//*****************************************************
// Project		: Fundamentals of class 1
// File			: section5_ex1_class1
// Editor		: Wenmei Wang
// Date			: 03/10/2024
// Description	: Fundamentals of class 1
//*****************************************************

class first;

	bit	[2:0]	data1;
	bit	[1:0]	data2;

endclass

module tb;

	first f;
	
	f.data1;
	f.data2;
	
endmodule