//*****************************************************
// Project		: Assignment 3 - A32
// File			: section3_a32
// Editor		: Wenmei Wang
// Date			: 21/09/2024
// Description	: Assignment 3 - A32
//*****************************************************

module tb;

	int arr[10] = '{0, 1, 4, 9, 16, 25, 36, 49, 64, 81};
	
	initial begin
		$display("arr : %0p", arr);
	end

endmodule