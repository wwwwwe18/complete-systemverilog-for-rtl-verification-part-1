//*****************************************************
// Project		: Injecting error
// File			: section8_ex7_inject_error
// Editor		: Wenmei Wang
// Date			: 13/10/2024
// Description	: Injecting error
//*****************************************************

class transaction;

	randc	bit	[3:0]	a;
	randc	bit	[3:0]	b;
			bit	[4:0]	sum;

	function void display();

		$display("a : %0d \t b : %0d \t sum : %0d", a, b, sum);

	endfunction

	virtual function transaction copy();	// Deep copy

		copy = new();
		copy.a = this.a;
		copy.b = this.b;
		copy.sum = this.sum;

	endfunction

endclass

class error extends transaction;

	//constraint	data_c	{a == 0; b == 0;}
	
	function transaction copy();

		copy = new();
		copy.a = 0;
		copy.b = 0;
		copy.sum = this.sum;

	endfunction

endclass

class generator;

	transaction trans;
	mailbox #(transaction) mbx;

	event done;

	int i = 0;

	function new(mailbox #(transaction) mbx);

		this.mbx = mbx;
		trans = new();

	endfunction

	task run();

		for(i = 0; i < 10; i++) begin

			trans.randomize();
			mbx.put(trans.copy);
			$display("[GEN] : DATA SENT TO DRIVER");
			trans.display();
			#20;

		end

		-> done;

	endtask

endclass

interface add_if;

	logic	[3:0]	a;
	logic	[3:0]	b;
	logic	[4:0]	sum;
	logic			clk;

endinterface

class driver;

	virtual add_if aif;	// Access interface
	mailbox #(transaction) mbx;
	transaction dc;
	event next;

	function new(mailbox #(transaction) mbx);

		this.mbx = mbx;

	endfunction

	task run();

		forever begin

			mbx.get(dc);
			@(posedge aif.clk);
			aif.a <= dc.a;
			aif.b <= dc.b;
			$display("[DRV] : Interface Trigger");
			dc.display();

		end

	endtask

endclass

module tb;

	add_if aif();
	driver drv;
	generator gen;
	error err;

	event done;

	mailbox #(transaction) mbx;

	add dut (.b(aif.b), .a(aif.a), .sum(aif.sum), .clk(aif.clk));

	initial begin

		aif.clk <= 0;

	end

	always #10 aif.clk <= ~aif.clk;

	initial begin

		mbx = new();
		err = new();
		gen = new(mbx);
		
		gen.trans = err;
		
		drv = new(mbx);
		drv.aif = aif;	// Connect interface in class to interface in tb
		done = gen.done;
		
	end

	initial begin

		fork

			gen.run();
			drv.run();

		join_none

		wait(done.triggered);
		$finish();

	end

	initial begin

		$dumpfile("dump.vcd");
		$dumpvars;

	end

endmodule