//*****************************************************
// Project		: Queue 1
// File			: section3_ex19_queue1
// Editor		: Wenmei Wang
// Date			: 01/10/2024
// Description	: Queue 1
//*****************************************************

module tb;

	int arr[$];
	
	initial begin
		arr = {1,2,3};
		$display("arr : %0p", arr);
	end

endmodule